module ctrl_unit (
    
);
    
endmodule